.subckt kicad_builtin_vdiff in+ in- out
  Emeas out 0 in+ in- 1
.ends